 `define no_of_trans 20
